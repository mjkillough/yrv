module yrv_top(
	input  [17:0] SW,
	output [17:0] LEDR
	);

    wire clk;
    wire res;

endmodule
